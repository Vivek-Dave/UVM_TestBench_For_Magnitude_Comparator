
interface intf();
    // ------------------- port declaration-------------------------------------
    logic [7:0] a;
    logic [7:0] b;
    logic     aeb;
    logic     alb;
    logic     agb;
    logic    aleb;
    logic    ageb;
    logic    aneb;
    //--------------------------------------------------------------------------
        
endinterface

