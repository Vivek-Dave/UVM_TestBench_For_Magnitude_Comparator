
`include "interface.sv"
`include "tb_pkg.sv"
module top;
  import uvm_pkg::*;
  import tb_pkg::*;
  
  //----------------------------------------------------------------------------
  intf i_intf();
  //----------------------------------------------------------------------------

  //----------------------------------------------------------------------------
  comparator DUT(.a(i_intf.a),
                 .b(i_intf.b),
                 .aeb(i_intf.aeb),
                 .alb(i_intf.alb),
                 .agb(i_intf.agb),
                 .aneb(i_intf.aneb),
                 .aleb(i_intf.aleb),
                 .ageb(i_intf.ageb)
                );
  //----------------------------------------------------------------------------               
  
  //----------------------------------------------------------------------------
  initial begin
    $dumpfile("dumpfile.vcd");
    $dumpvars;
  end
  //----------------------------------------------------------------------------

  //----------------------------------------------------------------------------
  initial begin
    uvm_config_db#(virtual intf)::set(uvm_root::get(),"","vif",i_intf);
  end
  //----------------------------------------------------------------------------

  //----------------------------------------------------------------------------
  initial begin
    run_test("comparator_test");
  end
  //----------------------------------------------------------------------------
endmodule

